module inv(y, x);
  (* src = "inverter/inverter.v:1.27-1.28" *)
  input x;
  wire x;
  (* src = "inverter/inverter.v:1.19-1.20" *)
  output y;
  wire y;
  INV_X1 _0_ (
    .A(x),
    .ZN(y)
  );
endmodule
