module inv(output y,input x);
not g1(y,x);
endmodule
